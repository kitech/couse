module mgs

fn test_build() {
	// println(sizeof(mg_mgr))
}
