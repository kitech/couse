module mongoose

fn test_build() {
	// println(sizeof(mg_mgr))
}
